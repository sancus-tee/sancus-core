module alias(.a(x), .b(x));
inout x;
wire x;
endmodule

